/**
 * ============================================================================
 * 寄存器堆模块 (Register File)
 * ============================================================================
 * 功能：
 * - 提供 32 个 32-bit 通用寄存器 (x0-x31)
 * - x0 固定为 0 (硬编码为零寄存器)
 * - 支持双端口读取 (Rs1, Rs2)
 * - 支持单端口写入 (Rd)
 * - 写优先读：同周期写入的数据可在同周期读出
 *
 * RISC-V 规范：
 * - x0 始终读为 0，写入 x0 无效
 * - 其他寄存器 x1-x31 可读可写
 * ============================================================================
 */

module regfile
    import rv32i_types::*;
    (
        input  logic        clk,        // 时钟信号
        input  logic        rst,        // 复位信号

        // ====================================================================
        // 写入接口 (来自 CDB)
        // ====================================================================
        input  logic        regf_we,    // 写使能
        input  logic [31:0] rd_v,       // 写入数据
        input  logic [4:0]  rd_s,       // 写入寄存器地址

        // ====================================================================
        // 读取接口 (到 Scoreboard)
        // ====================================================================
        input  logic [4:0]  rs1_s,      // Rs1 地址
        input  logic [4:0]  rs2_s,      // Rs2 地址
        output logic [31:0] rs1_v,      // Rs1 数据
        output logic [31:0] rs2_v       // Rs2 数据
    );

    // ========================================================================
    // 寄存器存储阵列
    // ========================================================================
    logic [31:0] data [32];

    // ========================================================================
    // 寄存器写入逻辑 (时序逻辑)
    // ========================================================================
    always_ff @(posedge clk) begin
        if (rst) begin
            // ----------------------------------------------------------------
            // 复位：清空所有寄存器
            // ----------------------------------------------------------------
            for (int i = 0; i < 32; i++) begin
                data[i] <= 32'b0;
            end

        end else if (regf_we && (rd_s != 5'd0)) begin
            // ----------------------------------------------------------------
            // 写入：只有 Rd 不是 x0 且写使能有效时才写入
            // ----------------------------------------------------------------
            data[rd_s] <= rd_v;
        end
    end

    // ========================================================================
    // 寄存器读取逻辑 (组合逻辑 + 写优先读)
    // ========================================================================
    always_comb begin
        // ----------------------------------------------------------------
        // Rs1 读取
        // ----------------------------------------------------------------
        if (rs1_s == 5'd0) begin
            // x0 寄存器始终为 0
            rs1_v = 32'b0;
        end else if (regf_we && (rs1_s == rd_s)) begin
            // 写优先读：同周期写入的数据直接转发
            rs1_v = rd_v;
        end else begin
            // 正常读取
            rs1_v = data[rs1_s];
        end

        // ----------------------------------------------------------------
        // Rs2 读取
        // ----------------------------------------------------------------
        if (rs2_s == 5'd0) begin
            rs2_v = 32'b0;
        end else if (regf_we && (rs2_s == rd_s)) begin
            rs2_v = rd_v;
        end else begin
            rs2_v = data[rs2_s];
        end
    end

endmodule : regfile
