/**
 * ============================================================================
 * 取指令阶段 (Fetch Stage)
 * ============================================================================
 * 功能：
 * - 从指令内存取指令
 * - 维护程序计数器 (PC)
 * - 处理分支跳转
 * - 将指令推入指令队列
 *
 * 控制流：
 * - 正常情况：PC = PC + 4
 * - 分支跳转：PC = branch_target (来自 Branch FU)
 * - 队列满：停止取指令 (反压)
 * ============================================================================
 */

module fetch
    import rv32i_types::*;
    (
        input  logic        clk,
        input  logic        rst,

        // ====================================================================
        // 指令内存接口
        // ====================================================================
        output logic [31:0] imem_addr,      // 取指地址
        output logic [3:0]  imem_rmask,     // 读掩码 (始终为 4'b1111)
        input  logic [31:0] imem_rdata,     // 指令数据
        input  logic        imem_resp,      // 内存响应

        // ====================================================================
        // 分支跳转接口 (来自 Branch FU)
        // ====================================================================
        input  logic        branch_taken,   // 分支是否跳转
        input  logic [31:0] branch_target,  // 分支目标地址

        // ====================================================================
        // 指令队列接口
        // ====================================================================
        output logic        iq_enq,         // 入队使能
        output iq_entry_t   iq_enq_data,    // 入队数据
        input  logic        iq_full         // 队列满标志
    );

    // ========================================================================
    // 程序计数器 (PC)
    // ========================================================================
    logic [31:0] pc, next_pc;

    // PC 初始值：RISC-V 规范要求从 0x60000000 开始
    localparam logic [31:0] PC_RESET_VALUE = 32'h60000000;

    always_ff @(posedge clk) begin
        if (rst) begin
            pc <= PC_RESET_VALUE;
        end else if (!iq_full && imem_resp) begin
            // 只有队列不满且内存响应时才更新 PC
            pc <= next_pc;
        end
    end

    // ========================================================================
    // 下一个 PC 计算 (组合逻辑)
    // ========================================================================
    always_comb begin
        if (branch_taken) begin
            // 分支跳转：跳转到目标地址
            next_pc = branch_target;
        end else begin
            // 正常情况：PC + 4
            next_pc = pc + 4;
        end
    end

    // ========================================================================
    // 指令内存访问
    // ========================================================================
    assign imem_addr = pc;
    assign imem_rmask = 4'b1111;  // 始终读取完整的 32-bit 字

    // ========================================================================
    // 指令序号追踪 (用于 RVFI 验证)
    // ========================================================================
    logic [63:0] instruction_order;

    always_ff @(posedge clk) begin
        if (rst) begin
            instruction_order <= 64'b0;
        end else if (iq_enq) begin
            instruction_order <= instruction_order + 1;
        end
    end

    // ========================================================================
    // 指令队列入队逻辑
    // ========================================================================
    assign iq_enq = imem_resp && !iq_full;

    always_comb begin
        iq_enq_data.inst  = imem_rdata;
        iq_enq_data.pc    = pc;
        iq_enq_data.order = instruction_order;
        iq_enq_data.valid = 1'b1;
    end

endmodule : fetch
